`include "const_arith_wrapper.sv"
`include "const_compare_wrapper.sv"
`include "const_concat_repl_wrapper.sv"
`include "const_conditional_wrapper.sv"
`include "const_logic_wrapper.sv"
`include "const_nested_wrapper.sv"
`include "const_partselect_wrapper.sv"
`include "const_reduce_wrapper.sv"
`include "const_shift_wrapper.sv"
`include "numbers_arithmetic_reduce_wrapper.sv"
`include "numbers_bitwise_logic_wrapper.sv"
`include "numbers_bitwise_reduce_wrapper.sv"
`include "numbers_concat_repl_wrapper.sv"
`include "numbers_constant_wrapper.sv"
`include "numbers_logical_op_wrapper.sv"
`include "numbers_numbers_arithmetic_wrapper.sv"
`include "numbers_reduce_case_wrapper.sv"
`include "numbers_relational_wrapper.sv"
`include "numbers_select_wrapper.sv"
`include "numbers_shift_wrapper.sv"
`include "widths_arith_wrapper.sv"
`include "widths_array_wrapper.sv"
`include "widths_cast_wrapper.sv"
`include "widths_concat_repl_wrapper.sv"
`include "widths_conditional_wrapper.sv"
`include "widths_enum_mod_wrapper.sv"
`include "widths_logic_mod_wrapper.sv"
`include "widths_param_wrapper.sv"
`include "widths_partselect_wrapper.sv"
`include "widths_shift_wrapper.sv"
`include "widths_struct_mod_wrapper.sv"
`include "widths_union_mod_wrapper.sv"

// Automatically generated top module
module top (
    input  wire [4:0] in_flat,
    output wire [476:0] out_flat
);

  // Per-module flattened I/O buses
  wire [15:0] const_arith_wrapper_in_flat;
  wire [39:0] const_arith_wrapper_out_flat;
  wire [23:0] const_compare_wrapper_in_flat;
  wire [7:0] const_compare_wrapper_out_flat;
  wire [9:0] const_concat_repl_wrapper_in_flat;
  wire [21:0] const_concat_repl_wrapper_out_flat;
  wire [33:0] const_conditional_wrapper_in_flat;
  wire [23:0] const_conditional_wrapper_out_flat;
  wire [9:0] const_logic_wrapper_in_flat;
  wire [18:0] const_logic_wrapper_out_flat;
  wire [26:0] const_nested_wrapper_in_flat;
  wire [7:0] const_nested_wrapper_out_flat;
  wire [19:0] const_partselect_wrapper_in_flat;
  wire [7:0] const_partselect_wrapper_out_flat;
  wire [3:0] const_reduce_wrapper_in_flat;
  wire [5:0] const_reduce_wrapper_out_flat;
  wire [10:0] const_shift_wrapper_in_flat;
  wire [23:0] const_shift_wrapper_out_flat;
  wire [15:0] numbers_arithmetic_reduce_wrapper_in_flat;
  wire [9:0] numbers_arithmetic_reduce_wrapper_out_flat;
  wire [15:0] numbers_bitwise_logic_wrapper_in_flat;
  wire [23:0] numbers_bitwise_logic_wrapper_out_flat;
  wire [7:0] numbers_bitwise_reduce_wrapper_in_flat;
  wire [2:0] numbers_bitwise_reduce_wrapper_out_flat;
  wire [5:0] numbers_concat_repl_wrapper_in_flat;
  wire [21:0] numbers_concat_repl_wrapper_out_flat;
  wire [0:0] numbers_constant_wrapper_in_flat;
  wire [79:0] numbers_constant_wrapper_out_flat;
  wire [1:0] numbers_logical_op_wrapper_in_flat;
  wire [2:0] numbers_logical_op_wrapper_out_flat;
  wire [12:0] numbers_numbers_arithmetic_wrapper_in_flat;
  wire [24:0] numbers_numbers_arithmetic_wrapper_out_flat;
  wire [7:0] numbers_reduce_case_wrapper_in_flat;
  wire [1:0] numbers_reduce_case_wrapper_out_flat;
  wire [7:0] numbers_relational_wrapper_in_flat;
  wire [7:0] numbers_relational_wrapper_out_flat;
  wire [19:0] numbers_select_wrapper_in_flat;
  wire [8:0] numbers_select_wrapper_out_flat;
  wire [10:0] numbers_shift_wrapper_in_flat;
  wire [15:0] numbers_shift_wrapper_out_flat;
  wire [0:0] widths_arith_wrapper_in_flat;
  wire [0:0] widths_arith_wrapper_out_flat;
  wire [17:0] widths_array_wrapper_in_flat;
  wire [15:0] widths_array_wrapper_out_flat;
  wire [11:0] widths_cast_wrapper_in_flat;
  wire [11:0] widths_cast_wrapper_out_flat;
  wire [5:0] widths_concat_repl_wrapper_in_flat;
  wire [17:0] widths_concat_repl_wrapper_out_flat;
  wire [8:0] widths_conditional_wrapper_in_flat;
  wire [3:0] widths_conditional_wrapper_out_flat;
  wire [3:0] widths_enum_mod_wrapper_in_flat;
  wire [4:0] widths_enum_mod_wrapper_out_flat;
  wire [7:0] widths_logic_mod_wrapper_in_flat;
  wire [5:0] widths_logic_mod_wrapper_out_flat;
  wire [0:0] widths_param_wrapper_in_flat;
  wire [0:0] widths_param_wrapper_out_flat;
  wire [18:0] widths_partselect_wrapper_in_flat;
  wire [8:0] widths_partselect_wrapper_out_flat;
  wire [10:0] widths_shift_wrapper_in_flat;
  wire [15:0] widths_shift_wrapper_out_flat;
  wire [11:0] widths_struct_mod_wrapper_in_flat;
  wire [11:0] widths_struct_mod_wrapper_out_flat;
  wire [15:0] widths_union_mod_wrapper_in_flat;
  wire [15:0] widths_union_mod_wrapper_out_flat;

  // Drive module inputs from top-level in_flat
  assign widths_struct_mod_wrapper_in_flat[4] = in_flat[2];
  assign numbers_bitwise_reduce_wrapper_in_flat[1] = in_flat[4];
  assign numbers_arithmetic_reduce_wrapper_in_flat[1] = in_flat[0];
  assign const_shift_wrapper_in_flat[6] = in_flat[3];
  assign const_reduce_wrapper_in_flat[1] = in_flat[1];

  // Internal connections: module-out → module-in
  assign widths_cast_wrapper_in_flat[4] = const_shift_wrapper_out_flat[15];
  assign widths_shift_wrapper_in_flat[0] = widths_cast_wrapper_out_flat[9];
  assign widths_struct_mod_wrapper_in_flat[1] = const_concat_repl_wrapper_out_flat[15];
  assign const_conditional_wrapper_in_flat[18] = const_logic_wrapper_out_flat[11];
  assign numbers_concat_repl_wrapper_in_flat[5] = const_shift_wrapper_out_flat[3];
  assign numbers_reduce_case_wrapper_in_flat[0] = numbers_arithmetic_reduce_wrapper_out_flat[8];
  assign const_arith_wrapper_in_flat[5] = widths_array_wrapper_out_flat[14];
  assign numbers_arithmetic_reduce_wrapper_in_flat[12] = const_reduce_wrapper_out_flat[1];
  assign numbers_numbers_arithmetic_wrapper_in_flat[10] = const_arith_wrapper_out_flat[25];
  assign const_partselect_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[15];
  assign const_nested_wrapper_in_flat[19] = widths_partselect_wrapper_out_flat[6];
  assign const_conditional_wrapper_in_flat[0] = widths_cast_wrapper_out_flat[1];
  assign widths_cast_wrapper_in_flat[9] = const_conditional_wrapper_out_flat[13];
  assign const_logic_wrapper_in_flat[6] = widths_shift_wrapper_out_flat[9];
  assign numbers_constant_wrapper_in_flat[0] = widths_concat_repl_wrapper_out_flat[0];
  assign const_conditional_wrapper_in_flat[14] = widths_shift_wrapper_out_flat[6];
  assign const_concat_repl_wrapper_in_flat[5] = numbers_constant_wrapper_out_flat[7];
  assign widths_enum_mod_wrapper_in_flat[2] = widths_logic_mod_wrapper_out_flat[0];
  assign widths_partselect_wrapper_in_flat[18] = numbers_numbers_arithmetic_wrapper_out_flat[7];
  assign numbers_select_wrapper_in_flat[13] = numbers_reduce_case_wrapper_out_flat[0];
  assign widths_partselect_wrapper_in_flat[16] = const_nested_wrapper_out_flat[5];
  assign const_partselect_wrapper_in_flat[10] = numbers_constant_wrapper_out_flat[45];
  assign widths_enum_mod_wrapper_in_flat[0] = numbers_constant_wrapper_out_flat[31];
  assign widths_partselect_wrapper_in_flat[1] = widths_partselect_wrapper_out_flat[2];
  assign const_concat_repl_wrapper_in_flat[8] = const_partselect_wrapper_out_flat[4];
  assign widths_logic_mod_wrapper_in_flat[2] = numbers_constant_wrapper_out_flat[19];
  assign const_arith_wrapper_in_flat[11] = numbers_arithmetic_reduce_wrapper_out_flat[4];
  assign numbers_bitwise_reduce_wrapper_in_flat[3] = const_concat_repl_wrapper_out_flat[9];
  assign numbers_bitwise_logic_wrapper_in_flat[11] = numbers_constant_wrapper_out_flat[42];
  assign numbers_numbers_arithmetic_wrapper_in_flat[4] = widths_enum_mod_wrapper_out_flat[0];
  assign const_conditional_wrapper_in_flat[12] = const_logic_wrapper_out_flat[17];
  assign widths_array_wrapper_in_flat[15] = const_concat_repl_wrapper_out_flat[6];
  assign numbers_bitwise_logic_wrapper_in_flat[5] = widths_struct_mod_wrapper_out_flat[2];
  assign numbers_concat_repl_wrapper_in_flat[2] = widths_cast_wrapper_out_flat[8];
  assign numbers_relational_wrapper_in_flat[4] = const_arith_wrapper_out_flat[37];
  assign numbers_select_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[16];
  assign widths_array_wrapper_in_flat[5] = const_compare_wrapper_out_flat[0];
  assign widths_shift_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[49];
  assign const_nested_wrapper_in_flat[14] = numbers_bitwise_reduce_wrapper_out_flat[1];
  assign widths_conditional_wrapper_in_flat[5] = const_logic_wrapper_out_flat[18];
  assign numbers_select_wrapper_in_flat[10] = const_logic_wrapper_out_flat[3];
  assign const_compare_wrapper_in_flat[5] = const_conditional_wrapper_out_flat[18];
  assign const_conditional_wrapper_in_flat[5] = widths_union_mod_wrapper_out_flat[5];
  assign numbers_numbers_arithmetic_wrapper_in_flat[5] = numbers_constant_wrapper_out_flat[64];
  assign widths_cast_wrapper_in_flat[1] = numbers_numbers_arithmetic_wrapper_out_flat[23];
  assign widths_partselect_wrapper_in_flat[10] = widths_partselect_wrapper_out_flat[5];
  assign const_partselect_wrapper_in_flat[12] = const_nested_wrapper_out_flat[7];
  assign const_compare_wrapper_in_flat[23] = numbers_constant_wrapper_out_flat[32];
  assign numbers_arithmetic_reduce_wrapper_in_flat[4] = const_concat_repl_wrapper_out_flat[1];
  assign widths_array_wrapper_in_flat[17] = numbers_constant_wrapper_out_flat[11];
  assign const_logic_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[27];
  assign numbers_bitwise_reduce_wrapper_in_flat[4] = widths_cast_wrapper_out_flat[11];
  assign widths_shift_wrapper_in_flat[2] = numbers_constant_wrapper_out_flat[0];
  assign numbers_bitwise_logic_wrapper_in_flat[13] = numbers_constant_wrapper_out_flat[57];
  assign const_partselect_wrapper_in_flat[9] = const_arith_wrapper_out_flat[15];
  assign numbers_numbers_arithmetic_wrapper_in_flat[1] = numbers_arithmetic_reduce_wrapper_out_flat[2];
  assign numbers_bitwise_reduce_wrapper_in_flat[0] = numbers_reduce_case_wrapper_out_flat[1];
  assign const_nested_wrapper_in_flat[7] = const_concat_repl_wrapper_out_flat[13];
  assign widths_cast_wrapper_in_flat[11] = const_arith_wrapper_out_flat[1];
  assign widths_cast_wrapper_in_flat[0] = const_partselect_wrapper_out_flat[1];
  assign const_partselect_wrapper_in_flat[3] = numbers_constant_wrapper_out_flat[56];
  assign widths_shift_wrapper_in_flat[10] = widths_array_wrapper_out_flat[4];
  assign const_compare_wrapper_in_flat[11] = widths_union_mod_wrapper_out_flat[12];
  assign numbers_arithmetic_reduce_wrapper_in_flat[9] = numbers_constant_wrapper_out_flat[51];
  assign const_compare_wrapper_in_flat[10] = numbers_concat_repl_wrapper_out_flat[15];
  assign const_partselect_wrapper_in_flat[19] = numbers_numbers_arithmetic_wrapper_out_flat[24];
  assign widths_concat_repl_wrapper_in_flat[5] = widths_struct_mod_wrapper_out_flat[0];
  assign const_partselect_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[8];
  assign const_nested_wrapper_in_flat[11] = numbers_concat_repl_wrapper_out_flat[19];
  assign widths_partselect_wrapper_in_flat[8] = const_arith_wrapper_out_flat[8];
  assign numbers_bitwise_logic_wrapper_in_flat[1] = numbers_numbers_arithmetic_wrapper_out_flat[22];
  assign const_partselect_wrapper_in_flat[18] = numbers_constant_wrapper_out_flat[34];
  assign numbers_numbers_arithmetic_wrapper_in_flat[2] = widths_conditional_wrapper_out_flat[1];
  assign const_shift_wrapper_in_flat[0] = const_conditional_wrapper_out_flat[7];
  assign const_partselect_wrapper_in_flat[14] = widths_param_wrapper_out_flat[0];
  assign numbers_reduce_case_wrapper_in_flat[1] = numbers_select_wrapper_out_flat[0];
  assign widths_array_wrapper_in_flat[8] = numbers_constant_wrapper_out_flat[70];
  assign numbers_arithmetic_reduce_wrapper_in_flat[3] = widths_struct_mod_wrapper_out_flat[5];
  assign const_compare_wrapper_in_flat[13] = const_arith_wrapper_out_flat[20];
  assign numbers_select_wrapper_in_flat[8] = numbers_shift_wrapper_out_flat[4];
  assign widths_union_mod_wrapper_in_flat[15] = numbers_bitwise_logic_wrapper_out_flat[5];
  assign widths_struct_mod_wrapper_in_flat[8] = widths_union_mod_wrapper_out_flat[8];
  assign const_concat_repl_wrapper_in_flat[4] = numbers_constant_wrapper_out_flat[76];
  assign numbers_shift_wrapper_in_flat[6] = numbers_relational_wrapper_out_flat[3];
  assign numbers_concat_repl_wrapper_in_flat[3] = const_arith_wrapper_out_flat[28];
  assign const_compare_wrapper_in_flat[6] = const_arith_wrapper_out_flat[6];
  assign numbers_numbers_arithmetic_wrapper_in_flat[3] = widths_array_wrapper_out_flat[15];
  assign widths_logic_mod_wrapper_in_flat[6] = numbers_numbers_arithmetic_wrapper_out_flat[1];
  assign numbers_relational_wrapper_in_flat[2] = numbers_shift_wrapper_out_flat[12];
  assign widths_partselect_wrapper_in_flat[17] = widths_shift_wrapper_out_flat[11];
  assign const_compare_wrapper_in_flat[7] = const_conditional_wrapper_out_flat[11];
  assign const_arith_wrapper_in_flat[4] = numbers_constant_wrapper_out_flat[60];
  assign const_conditional_wrapper_in_flat[6] = numbers_select_wrapper_out_flat[8];
  assign numbers_concat_repl_wrapper_in_flat[0] = const_arith_wrapper_out_flat[39];
  assign const_partselect_wrapper_in_flat[6] = numbers_arithmetic_reduce_wrapper_out_flat[0];
  assign const_nested_wrapper_in_flat[8] = widths_shift_wrapper_out_flat[7];
  assign const_nested_wrapper_in_flat[2] = numbers_bitwise_logic_wrapper_out_flat[9];
  assign const_conditional_wrapper_in_flat[25] = numbers_numbers_arithmetic_wrapper_out_flat[11];
  assign numbers_select_wrapper_in_flat[19] = const_conditional_wrapper_out_flat[15];
  assign const_nested_wrapper_in_flat[5] = const_conditional_wrapper_out_flat[6];
  assign widths_logic_mod_wrapper_in_flat[0] = const_conditional_wrapper_out_flat[19];
  assign numbers_arithmetic_reduce_wrapper_in_flat[0] = widths_union_mod_wrapper_out_flat[15];
  assign const_nested_wrapper_in_flat[22] = widths_logic_mod_wrapper_out_flat[3];
  assign widths_cast_wrapper_in_flat[7] = widths_union_mod_wrapper_out_flat[11];
  assign widths_enum_mod_wrapper_in_flat[3] = widths_concat_repl_wrapper_out_flat[15];
  assign widths_union_mod_wrapper_in_flat[12] = widths_union_mod_wrapper_out_flat[10];
  assign widths_union_mod_wrapper_in_flat[1] = widths_struct_mod_wrapper_out_flat[8];
  assign numbers_bitwise_reduce_wrapper_in_flat[2] = numbers_constant_wrapper_out_flat[43];
  assign const_nested_wrapper_in_flat[4] = const_shift_wrapper_out_flat[10];
  assign widths_struct_mod_wrapper_in_flat[11] = widths_cast_wrapper_out_flat[0];
  assign const_shift_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[72];
  assign const_conditional_wrapper_in_flat[28] = widths_array_wrapper_out_flat[2];
  assign widths_arith_wrapper_in_flat[0] = const_compare_wrapper_out_flat[5];
  assign numbers_select_wrapper_in_flat[0] = numbers_shift_wrapper_out_flat[9];
  assign widths_shift_wrapper_in_flat[3] = widths_union_mod_wrapper_out_flat[0];
  assign numbers_select_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[37];
  assign widths_struct_mod_wrapper_in_flat[6] = numbers_bitwise_logic_wrapper_out_flat[23];
  assign widths_union_mod_wrapper_in_flat[11] = const_conditional_wrapper_out_flat[20];
  assign numbers_numbers_arithmetic_wrapper_in_flat[12] = const_arith_wrapper_out_flat[38];
  assign numbers_bitwise_logic_wrapper_in_flat[12] = numbers_constant_wrapper_out_flat[47];
  assign numbers_arithmetic_reduce_wrapper_in_flat[13] = numbers_bitwise_logic_wrapper_out_flat[11];
  assign const_nested_wrapper_in_flat[9] = const_logic_wrapper_out_flat[16];
  assign const_concat_repl_wrapper_in_flat[0] = widths_array_wrapper_out_flat[5];
  assign const_conditional_wrapper_in_flat[21] = widths_shift_wrapper_out_flat[3];
  assign const_partselect_wrapper_in_flat[17] = numbers_relational_wrapper_out_flat[5];
  assign widths_cast_wrapper_in_flat[8] = const_arith_wrapper_out_flat[17];
  assign widths_union_mod_wrapper_in_flat[3] = const_logic_wrapper_out_flat[4];
  assign numbers_numbers_arithmetic_wrapper_in_flat[7] = numbers_arithmetic_reduce_wrapper_out_flat[1];
  assign const_arith_wrapper_in_flat[12] = numbers_numbers_arithmetic_wrapper_out_flat[20];
  assign widths_partselect_wrapper_in_flat[0] = const_logic_wrapper_out_flat[7];
  assign numbers_bitwise_logic_wrapper_in_flat[8] = const_logic_wrapper_out_flat[0];
  assign numbers_bitwise_logic_wrapper_in_flat[7] = const_arith_wrapper_out_flat[10];
  assign numbers_arithmetic_reduce_wrapper_in_flat[10] = const_shift_wrapper_out_flat[21];
  assign widths_concat_repl_wrapper_in_flat[0] = numbers_concat_repl_wrapper_out_flat[12];
  assign widths_shift_wrapper_in_flat[1] = widths_partselect_wrapper_out_flat[0];
  assign widths_cast_wrapper_in_flat[3] = numbers_bitwise_logic_wrapper_out_flat[8];
  assign numbers_select_wrapper_in_flat[6] = numbers_numbers_arithmetic_wrapper_out_flat[17];
  assign const_arith_wrapper_in_flat[14] = const_shift_wrapper_out_flat[13];
  assign widths_union_mod_wrapper_in_flat[4] = const_shift_wrapper_out_flat[19];
  assign const_arith_wrapper_in_flat[10] = numbers_bitwise_logic_wrapper_out_flat[15];
  assign numbers_bitwise_logic_wrapper_in_flat[4] = widths_cast_wrapper_out_flat[7];
  assign widths_logic_mod_wrapper_in_flat[3] = const_logic_wrapper_out_flat[2];
  assign const_arith_wrapper_in_flat[3] = numbers_bitwise_logic_wrapper_out_flat[10];
  assign widths_array_wrapper_in_flat[12] = const_arith_wrapper_out_flat[21];
  assign numbers_select_wrapper_in_flat[18] = widths_logic_mod_wrapper_out_flat[4];
  assign numbers_select_wrapper_in_flat[11] = const_concat_repl_wrapper_out_flat[0];
  assign const_nested_wrapper_in_flat[26] = const_nested_wrapper_out_flat[3];
  assign const_nested_wrapper_in_flat[6] = const_shift_wrapper_out_flat[2];
  assign const_partselect_wrapper_in_flat[0] = widths_logic_mod_wrapper_out_flat[2];
  assign const_conditional_wrapper_in_flat[13] = widths_union_mod_wrapper_out_flat[2];
  assign widths_union_mod_wrapper_in_flat[13] = numbers_constant_wrapper_out_flat[40];
  assign widths_partselect_wrapper_in_flat[11] = widths_concat_repl_wrapper_out_flat[12];
  assign const_compare_wrapper_in_flat[4] = numbers_concat_repl_wrapper_out_flat[21];
  assign const_partselect_wrapper_in_flat[2] = const_compare_wrapper_out_flat[4];
  assign widths_concat_repl_wrapper_in_flat[1] = widths_array_wrapper_out_flat[12];
  assign numbers_select_wrapper_in_flat[14] = const_compare_wrapper_out_flat[7];
  assign widths_array_wrapper_in_flat[3] = widths_partselect_wrapper_out_flat[8];
  assign const_nested_wrapper_in_flat[16] = widths_shift_wrapper_out_flat[10];
  assign const_arith_wrapper_in_flat[8] = const_shift_wrapper_out_flat[14];
  assign numbers_bitwise_logic_wrapper_in_flat[15] = numbers_constant_wrapper_out_flat[14];
  assign widths_struct_mod_wrapper_in_flat[0] = widths_array_wrapper_out_flat[9];
  assign numbers_shift_wrapper_in_flat[9] = widths_array_wrapper_out_flat[10];
  assign const_nested_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[20];
  assign widths_conditional_wrapper_in_flat[6] = numbers_constant_wrapper_out_flat[26];
  assign const_arith_wrapper_in_flat[13] = const_conditional_wrapper_out_flat[5];
  assign numbers_numbers_arithmetic_wrapper_in_flat[9] = numbers_constant_wrapper_out_flat[48];
  assign numbers_arithmetic_reduce_wrapper_in_flat[14] = numbers_concat_repl_wrapper_out_flat[13];
  assign const_arith_wrapper_in_flat[0] = widths_concat_repl_wrapper_out_flat[16];
  assign const_conditional_wrapper_in_flat[16] = numbers_constant_wrapper_out_flat[28];
  assign widths_union_mod_wrapper_in_flat[8] = widths_partselect_wrapper_out_flat[3];
  assign const_nested_wrapper_in_flat[21] = numbers_constant_wrapper_out_flat[46];
  assign numbers_relational_wrapper_in_flat[0] = const_concat_repl_wrapper_out_flat[21];
  assign widths_conditional_wrapper_in_flat[2] = const_logic_wrapper_out_flat[13];
  assign numbers_shift_wrapper_in_flat[5] = numbers_constant_wrapper_out_flat[75];
  assign const_conditional_wrapper_in_flat[9] = const_shift_wrapper_out_flat[1];
  assign const_conditional_wrapper_in_flat[29] = const_conditional_wrapper_out_flat[2];
  assign const_conditional_wrapper_in_flat[24] = numbers_concat_repl_wrapper_out_flat[16];
  assign const_logic_wrapper_in_flat[9] = const_concat_repl_wrapper_out_flat[20];
  assign numbers_reduce_case_wrapper_in_flat[3] = numbers_bitwise_reduce_wrapper_out_flat[2];
  assign const_nested_wrapper_in_flat[20] = numbers_constant_wrapper_out_flat[30];
  assign const_arith_wrapper_in_flat[6] = numbers_bitwise_logic_wrapper_out_flat[19];
  assign numbers_shift_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[10];
  assign widths_cast_wrapper_in_flat[5] = widths_cast_wrapper_out_flat[4];
  assign widths_struct_mod_wrapper_in_flat[7] = numbers_bitwise_logic_wrapper_out_flat[1];
  assign numbers_select_wrapper_in_flat[9] = const_concat_repl_wrapper_out_flat[10];
  assign numbers_reduce_case_wrapper_in_flat[2] = numbers_numbers_arithmetic_wrapper_out_flat[5];
  assign widths_concat_repl_wrapper_in_flat[2] = const_logic_wrapper_out_flat[9];
  assign const_partselect_wrapper_in_flat[15] = numbers_select_wrapper_out_flat[7];
  assign const_conditional_wrapper_in_flat[3] = numbers_arithmetic_reduce_wrapper_out_flat[3];
  assign widths_array_wrapper_in_flat[6] = numbers_constant_wrapper_out_flat[52];
  assign widths_concat_repl_wrapper_in_flat[4] = const_shift_wrapper_out_flat[17];
  assign numbers_relational_wrapper_in_flat[6] = const_concat_repl_wrapper_out_flat[11];
  assign numbers_logical_op_wrapper_in_flat[1] = const_logic_wrapper_out_flat[1];
  assign numbers_numbers_arithmetic_wrapper_in_flat[11] = numbers_constant_wrapper_out_flat[66];
  assign const_compare_wrapper_in_flat[15] = const_partselect_wrapper_out_flat[2];
  assign const_arith_wrapper_in_flat[9] = numbers_arithmetic_reduce_wrapper_out_flat[6];
  assign widths_array_wrapper_in_flat[7] = const_arith_wrapper_out_flat[16];
  assign widths_partselect_wrapper_in_flat[14] = const_conditional_wrapper_out_flat[9];
  assign const_conditional_wrapper_in_flat[1] = numbers_concat_repl_wrapper_out_flat[18];
  assign const_conditional_wrapper_in_flat[20] = widths_union_mod_wrapper_out_flat[3];
  assign widths_union_mod_wrapper_in_flat[2] = widths_struct_mod_wrapper_out_flat[4];
  assign const_shift_wrapper_in_flat[4] = widths_concat_repl_wrapper_out_flat[17];
  assign const_logic_wrapper_in_flat[5] = numbers_shift_wrapper_out_flat[14];
  assign widths_array_wrapper_in_flat[0] = numbers_shift_wrapper_out_flat[6];
  assign const_logic_wrapper_in_flat[8] = const_shift_wrapper_out_flat[7];
  assign numbers_shift_wrapper_in_flat[10] = const_logic_wrapper_out_flat[8];
  assign widths_union_mod_wrapper_in_flat[9] = numbers_concat_repl_wrapper_out_flat[17];
  assign numbers_select_wrapper_in_flat[17] = const_conditional_wrapper_out_flat[23];
  assign const_conditional_wrapper_in_flat[15] = const_conditional_wrapper_out_flat[16];
  assign const_compare_wrapper_in_flat[19] = const_conditional_wrapper_out_flat[14];
  assign widths_array_wrapper_in_flat[10] = numbers_numbers_arithmetic_wrapper_out_flat[19];
  assign const_compare_wrapper_in_flat[17] = numbers_constant_wrapper_out_flat[12];
  assign numbers_arithmetic_reduce_wrapper_in_flat[5] = numbers_constant_wrapper_out_flat[1];
  assign const_compare_wrapper_in_flat[3] = numbers_constant_wrapper_out_flat[71];
  assign widths_logic_mod_wrapper_in_flat[7] = widths_shift_wrapper_out_flat[2];
  assign widths_struct_mod_wrapper_in_flat[10] = const_conditional_wrapper_out_flat[17];
  assign widths_shift_wrapper_in_flat[4] = numbers_logical_op_wrapper_out_flat[1];
  assign widths_partselect_wrapper_in_flat[5] = const_reduce_wrapper_out_flat[0];
  assign widths_partselect_wrapper_in_flat[13] = const_conditional_wrapper_out_flat[0];
  assign numbers_arithmetic_reduce_wrapper_in_flat[2] = const_partselect_wrapper_out_flat[3];
  assign const_conditional_wrapper_in_flat[23] = numbers_numbers_arithmetic_wrapper_out_flat[6];
  assign numbers_bitwise_reduce_wrapper_in_flat[5] = const_conditional_wrapper_out_flat[12];
  assign widths_array_wrapper_in_flat[16] = const_concat_repl_wrapper_out_flat[3];
  assign numbers_reduce_case_wrapper_in_flat[7] = numbers_numbers_arithmetic_wrapper_out_flat[14];
  assign numbers_relational_wrapper_in_flat[7] = widths_shift_wrapper_out_flat[12];
  assign const_conditional_wrapper_in_flat[31] = widths_enum_mod_wrapper_out_flat[4];
  assign widths_array_wrapper_in_flat[9] = const_conditional_wrapper_out_flat[3];
  assign const_partselect_wrapper_in_flat[11] = widths_cast_wrapper_out_flat[3];
  assign widths_logic_mod_wrapper_in_flat[4] = widths_partselect_wrapper_out_flat[7];
  assign widths_partselect_wrapper_in_flat[9] = const_shift_wrapper_out_flat[5];
  assign numbers_relational_wrapper_in_flat[1] = const_arith_wrapper_out_flat[23];
  assign widths_array_wrapper_in_flat[4] = widths_cast_wrapper_out_flat[10];
  assign const_nested_wrapper_in_flat[13] = numbers_select_wrapper_out_flat[5];
  assign const_arith_wrapper_in_flat[7] = numbers_bitwise_logic_wrapper_out_flat[16];
  assign const_reduce_wrapper_in_flat[2] = numbers_constant_wrapper_out_flat[39];
  assign const_conditional_wrapper_in_flat[22] = widths_conditional_wrapper_out_flat[0];
  assign numbers_arithmetic_reduce_wrapper_in_flat[11] = numbers_concat_repl_wrapper_out_flat[11];
  assign numbers_select_wrapper_in_flat[12] = numbers_numbers_arithmetic_wrapper_out_flat[16];
  assign const_partselect_wrapper_in_flat[4] = numbers_constant_wrapper_out_flat[74];
  assign const_conditional_wrapper_in_flat[4] = numbers_arithmetic_reduce_wrapper_out_flat[9];
  assign const_concat_repl_wrapper_in_flat[2] = const_concat_repl_wrapper_out_flat[12];
  assign const_compare_wrapper_in_flat[8] = const_concat_repl_wrapper_out_flat[8];
  assign const_conditional_wrapper_in_flat[10] = widths_struct_mod_wrapper_out_flat[9];
  assign widths_union_mod_wrapper_in_flat[5] = widths_cast_wrapper_out_flat[2];
  assign widths_struct_mod_wrapper_in_flat[2] = numbers_arithmetic_reduce_wrapper_out_flat[7];
  assign widths_partselect_wrapper_in_flat[15] = numbers_select_wrapper_out_flat[3];
  assign numbers_reduce_case_wrapper_in_flat[5] = widths_enum_mod_wrapper_out_flat[3];
  assign const_shift_wrapper_in_flat[3] = const_arith_wrapper_out_flat[26];
  assign const_compare_wrapper_in_flat[12] = const_shift_wrapper_out_flat[22];
  assign const_concat_repl_wrapper_in_flat[1] = widths_logic_mod_wrapper_out_flat[5];
  assign numbers_shift_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[63];
  assign const_concat_repl_wrapper_in_flat[9] = numbers_numbers_arithmetic_wrapper_out_flat[2];
  assign widths_conditional_wrapper_in_flat[3] = const_shift_wrapper_out_flat[8];
  assign const_conditional_wrapper_in_flat[32] = widths_array_wrapper_out_flat[3];
  assign const_compare_wrapper_in_flat[1] = const_arith_wrapper_out_flat[18];
  assign const_conditional_wrapper_in_flat[11] = const_reduce_wrapper_out_flat[5];
  assign const_logic_wrapper_in_flat[3] = const_arith_wrapper_out_flat[31];
  assign const_nested_wrapper_in_flat[17] = widths_shift_wrapper_out_flat[13];
  assign const_shift_wrapper_in_flat[2] = numbers_shift_wrapper_out_flat[0];
  assign numbers_bitwise_logic_wrapper_in_flat[9] = numbers_constant_wrapper_out_flat[58];
  assign widths_partselect_wrapper_in_flat[2] = const_conditional_wrapper_out_flat[4];
  assign numbers_arithmetic_reduce_wrapper_in_flat[7] = const_logic_wrapper_out_flat[14];
  assign widths_partselect_wrapper_in_flat[3] = widths_conditional_wrapper_out_flat[3];
  assign widths_logic_mod_wrapper_in_flat[5] = numbers_concat_repl_wrapper_out_flat[10];
  assign widths_partselect_wrapper_in_flat[12] = numbers_arithmetic_reduce_wrapper_out_flat[5];
  assign const_shift_wrapper_in_flat[10] = numbers_numbers_arithmetic_wrapper_out_flat[0];
  assign widths_partselect_wrapper_in_flat[7] = numbers_concat_repl_wrapper_out_flat[1];
  assign widths_cast_wrapper_in_flat[6] = const_arith_wrapper_out_flat[32];
  assign widths_param_wrapper_in_flat[0] = numbers_concat_repl_wrapper_out_flat[2];
  assign numbers_shift_wrapper_in_flat[3] = widths_shift_wrapper_out_flat[1];
  assign const_nested_wrapper_in_flat[18] = widths_shift_wrapper_out_flat[8];
  assign const_nested_wrapper_in_flat[0] = widths_concat_repl_wrapper_out_flat[9];
  assign const_nested_wrapper_in_flat[23] = widths_union_mod_wrapper_out_flat[6];
  assign numbers_reduce_case_wrapper_in_flat[6] = const_concat_repl_wrapper_out_flat[5];
  assign numbers_logical_op_wrapper_in_flat[0] = widths_union_mod_wrapper_out_flat[9];
  assign widths_union_mod_wrapper_in_flat[6] = const_arith_wrapper_out_flat[13];
  assign numbers_bitwise_logic_wrapper_in_flat[0] = numbers_numbers_arithmetic_wrapper_out_flat[12];
  assign numbers_shift_wrapper_in_flat[2] = widths_array_wrapper_out_flat[6];
  assign numbers_arithmetic_reduce_wrapper_in_flat[15] = const_nested_wrapper_out_flat[2];
  assign const_conditional_wrapper_in_flat[7] = const_shift_wrapper_out_flat[20];
  assign const_nested_wrapper_in_flat[15] = numbers_concat_repl_wrapper_out_flat[4];
  assign widths_shift_wrapper_in_flat[9] = widths_partselect_wrapper_out_flat[1];
  assign numbers_bitwise_reduce_wrapper_in_flat[6] = numbers_bitwise_logic_wrapper_out_flat[14];
  assign widths_partselect_wrapper_in_flat[4] = widths_concat_repl_wrapper_out_flat[2];
  assign widths_concat_repl_wrapper_in_flat[3] = widths_logic_mod_wrapper_out_flat[1];
  assign widths_conditional_wrapper_in_flat[4] = numbers_bitwise_logic_wrapper_out_flat[4];
  assign const_nested_wrapper_in_flat[12] = const_shift_wrapper_out_flat[11];
  assign const_compare_wrapper_in_flat[21] = const_shift_wrapper_out_flat[0];
  assign const_logic_wrapper_in_flat[4] = const_compare_wrapper_out_flat[3];
  assign widths_array_wrapper_in_flat[13] = numbers_shift_wrapper_out_flat[10];
  assign numbers_select_wrapper_in_flat[2] = numbers_constant_wrapper_out_flat[38];
  assign const_arith_wrapper_in_flat[15] = widths_conditional_wrapper_out_flat[2];
  assign const_concat_repl_wrapper_in_flat[6] = const_arith_wrapper_out_flat[2];
  assign widths_conditional_wrapper_in_flat[1] = widths_cast_wrapper_out_flat[5];
  assign const_nested_wrapper_in_flat[10] = const_conditional_wrapper_out_flat[21];
  assign const_compare_wrapper_in_flat[0] = numbers_shift_wrapper_out_flat[15];
  assign widths_struct_mod_wrapper_in_flat[9] = const_arith_wrapper_out_flat[11];
  assign const_logic_wrapper_in_flat[0] = widths_struct_mod_wrapper_out_flat[11];
  assign widths_union_mod_wrapper_in_flat[7] = numbers_constant_wrapper_out_flat[69];
  assign widths_array_wrapper_in_flat[1] = widths_union_mod_wrapper_out_flat[4];
  assign const_reduce_wrapper_in_flat[0] = const_shift_wrapper_out_flat[4];
  assign numbers_select_wrapper_in_flat[15] = numbers_relational_wrapper_out_flat[7];
  assign numbers_numbers_arithmetic_wrapper_in_flat[6] = numbers_bitwise_logic_wrapper_out_flat[3];
  assign widths_shift_wrapper_in_flat[8] = numbers_concat_repl_wrapper_out_flat[0];
  assign const_partselect_wrapper_in_flat[5] = numbers_logical_op_wrapper_out_flat[0];
  assign const_partselect_wrapper_in_flat[13] = widths_cast_wrapper_out_flat[6];
  assign numbers_select_wrapper_in_flat[3] = numbers_concat_repl_wrapper_out_flat[8];
  assign const_shift_wrapper_in_flat[1] = widths_union_mod_wrapper_out_flat[7];
  assign widths_union_mod_wrapper_in_flat[10] = numbers_constant_wrapper_out_flat[4];
  assign numbers_shift_wrapper_in_flat[0] = widths_struct_mod_wrapper_out_flat[1];
  assign const_partselect_wrapper_in_flat[16] = const_arith_wrapper_out_flat[9];
  assign numbers_select_wrapper_in_flat[5] = numbers_constant_wrapper_out_flat[21];
  assign const_compare_wrapper_in_flat[9] = numbers_constant_wrapper_out_flat[3];
  assign const_arith_wrapper_in_flat[1] = const_arith_wrapper_out_flat[7];
  assign numbers_relational_wrapper_in_flat[3] = const_logic_wrapper_out_flat[10];
  assign const_conditional_wrapper_in_flat[26] = numbers_shift_wrapper_out_flat[11];
  assign widths_union_mod_wrapper_in_flat[14] = numbers_constant_wrapper_out_flat[29];
  assign widths_partselect_wrapper_in_flat[6] = numbers_bitwise_logic_wrapper_out_flat[6];
  assign const_conditional_wrapper_in_flat[2] = widths_array_wrapper_out_flat[0];
  assign widths_conditional_wrapper_in_flat[8] = numbers_constant_wrapper_out_flat[35];
  assign numbers_numbers_arithmetic_wrapper_in_flat[0] = numbers_constant_wrapper_out_flat[41];
  assign const_reduce_wrapper_in_flat[3] = widths_shift_wrapper_out_flat[4];
  assign const_nested_wrapper_in_flat[25] = const_partselect_wrapper_out_flat[5];
  assign widths_array_wrapper_in_flat[2] = numbers_relational_wrapper_out_flat[0];
  assign const_conditional_wrapper_in_flat[27] = widths_array_wrapper_out_flat[8];
  assign const_conditional_wrapper_in_flat[17] = numbers_shift_wrapper_out_flat[8];
  assign widths_shift_wrapper_in_flat[6] = widths_array_wrapper_out_flat[13];
  assign numbers_reduce_case_wrapper_in_flat[4] = numbers_bitwise_logic_wrapper_out_flat[20];
  assign numbers_arithmetic_reduce_wrapper_in_flat[6] = numbers_numbers_arithmetic_wrapper_out_flat[8];
  assign const_concat_repl_wrapper_in_flat[7] = widths_enum_mod_wrapper_out_flat[2];
  assign const_nested_wrapper_in_flat[3] = numbers_constant_wrapper_out_flat[79];
  assign widths_struct_mod_wrapper_in_flat[3] = numbers_shift_wrapper_out_flat[5];
  assign numbers_concat_repl_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[13];
  assign const_concat_repl_wrapper_in_flat[3] = numbers_select_wrapper_out_flat[1];
  assign numbers_numbers_arithmetic_wrapper_in_flat[8] = numbers_bitwise_logic_wrapper_out_flat[18];
  assign const_conditional_wrapper_in_flat[19] = numbers_concat_repl_wrapper_out_flat[20];
  assign numbers_concat_repl_wrapper_in_flat[4] = numbers_numbers_arithmetic_wrapper_out_flat[15];
  assign const_partselect_wrapper_in_flat[8] = const_arith_wrapper_out_flat[22];
  assign widths_logic_mod_wrapper_in_flat[1] = numbers_constant_wrapper_out_flat[9];
  assign widths_conditional_wrapper_in_flat[7] = widths_concat_repl_wrapper_out_flat[13];
  assign numbers_select_wrapper_in_flat[16] = numbers_bitwise_reduce_wrapper_out_flat[0];
  assign const_nested_wrapper_in_flat[24] = widths_concat_repl_wrapper_out_flat[10];
  assign numbers_relational_wrapper_in_flat[5] = const_nested_wrapper_out_flat[1];
  assign numbers_bitwise_logic_wrapper_in_flat[14] = numbers_relational_wrapper_out_flat[2];
  assign const_logic_wrapper_in_flat[2] = widths_shift_wrapper_out_flat[0];
  assign numbers_bitwise_logic_wrapper_in_flat[6] = numbers_constant_wrapper_out_flat[77];
  assign const_compare_wrapper_in_flat[16] = numbers_constant_wrapper_out_flat[59];
  assign const_shift_wrapper_in_flat[8] = widths_union_mod_wrapper_out_flat[14];
  assign const_compare_wrapper_in_flat[20] = const_conditional_wrapper_out_flat[22];
  assign numbers_bitwise_logic_wrapper_in_flat[2] = widths_array_wrapper_out_flat[11];
  assign numbers_bitwise_logic_wrapper_in_flat[10] = numbers_constant_wrapper_out_flat[17];
  assign numbers_shift_wrapper_in_flat[4] = numbers_shift_wrapper_out_flat[3];
  assign widths_struct_mod_wrapper_in_flat[5] = widths_concat_repl_wrapper_out_flat[11];
  assign const_shift_wrapper_in_flat[9] = numbers_numbers_arithmetic_wrapper_out_flat[4];
  assign const_shift_wrapper_in_flat[5] = numbers_shift_wrapper_out_flat[2];
  assign const_conditional_wrapper_in_flat[30] = const_concat_repl_wrapper_out_flat[14];
  assign widths_cast_wrapper_in_flat[10] = const_partselect_wrapper_out_flat[6];
  assign widths_conditional_wrapper_in_flat[0] = const_arith_wrapper_out_flat[19];
  assign const_compare_wrapper_in_flat[14] = numbers_relational_wrapper_out_flat[6];
  assign numbers_bitwise_logic_wrapper_in_flat[3] = const_arith_wrapper_out_flat[33];
  assign widths_array_wrapper_in_flat[14] = widths_concat_repl_wrapper_out_flat[5];
  assign const_arith_wrapper_in_flat[2] = const_arith_wrapper_out_flat[3];
  assign widths_shift_wrapper_in_flat[5] = const_arith_wrapper_out_flat[4];
  assign numbers_shift_wrapper_in_flat[8] = numbers_constant_wrapper_out_flat[53];
  assign const_compare_wrapper_in_flat[22] = const_concat_repl_wrapper_out_flat[2];
  assign const_conditional_wrapper_in_flat[33] = numbers_constant_wrapper_out_flat[18];
  assign const_conditional_wrapper_in_flat[8] = numbers_constant_wrapper_out_flat[25];
  assign numbers_select_wrapper_in_flat[4] = numbers_constant_wrapper_out_flat[36];
  assign widths_cast_wrapper_in_flat[2] = const_compare_wrapper_out_flat[2];
  assign const_compare_wrapper_in_flat[18] = const_shift_wrapper_out_flat[18];
  assign numbers_arithmetic_reduce_wrapper_in_flat[8] = numbers_concat_repl_wrapper_out_flat[14];
  assign widths_union_mod_wrapper_in_flat[0] = numbers_bitwise_logic_wrapper_out_flat[12];
  assign numbers_bitwise_reduce_wrapper_in_flat[7] = const_logic_wrapper_out_flat[6];
  assign widths_array_wrapper_in_flat[11] = numbers_bitwise_logic_wrapper_out_flat[22];
  assign widths_enum_mod_wrapper_in_flat[1] = numbers_select_wrapper_out_flat[4];
  assign const_compare_wrapper_in_flat[2] = widths_enum_mod_wrapper_out_flat[1];
  assign const_logic_wrapper_in_flat[7] = widths_concat_repl_wrapper_out_flat[14];

  // Drive top-level out_flat from module outputs
  assign out_flat[423] = numbers_relational_wrapper_out_flat[0];
  assign out_flat[81] = numbers_relational_wrapper_out_flat[1];
  assign out_flat[443] = numbers_relational_wrapper_out_flat[2];
  assign out_flat[183] = numbers_relational_wrapper_out_flat[3];
  assign out_flat[66] = numbers_relational_wrapper_out_flat[4];
  assign out_flat[224] = numbers_relational_wrapper_out_flat[5];
  assign out_flat[458] = numbers_relational_wrapper_out_flat[6];
  assign out_flat[401] = numbers_relational_wrapper_out_flat[7];
  assign out_flat[403] = numbers_concat_repl_wrapper_out_flat[0];
  assign out_flat[366] = numbers_concat_repl_wrapper_out_flat[1];
  assign out_flat[368] = numbers_concat_repl_wrapper_out_flat[2];
  assign out_flat[70] = numbers_concat_repl_wrapper_out_flat[3];
  assign out_flat[380] = numbers_concat_repl_wrapper_out_flat[4];
  assign out_flat[69] = numbers_concat_repl_wrapper_out_flat[5];
  assign out_flat[89] = numbers_concat_repl_wrapper_out_flat[6];
  assign out_flat[71] = numbers_concat_repl_wrapper_out_flat[7];
  assign out_flat[406] = numbers_concat_repl_wrapper_out_flat[8];
  assign out_flat[19] = numbers_concat_repl_wrapper_out_flat[9];
  assign out_flat[363] = numbers_concat_repl_wrapper_out_flat[10];
  assign out_flat[336] = numbers_concat_repl_wrapper_out_flat[11];
  assign out_flat[233] = numbers_concat_repl_wrapper_out_flat[12];
  assign out_flat[266] = numbers_concat_repl_wrapper_out_flat[13];
  assign out_flat[470] = numbers_concat_repl_wrapper_out_flat[14];
  assign out_flat[164] = numbers_concat_repl_wrapper_out_flat[15];
  assign out_flat[276] = numbers_concat_repl_wrapper_out_flat[16];
  assign out_flat[306] = numbers_concat_repl_wrapper_out_flat[17];
  assign out_flat[298] = numbers_concat_repl_wrapper_out_flat[18];
  assign out_flat[168] = numbers_concat_repl_wrapper_out_flat[19];
  assign out_flat[435] = numbers_concat_repl_wrapper_out_flat[20];
  assign out_flat[252] = numbers_concat_repl_wrapper_out_flat[21];
  assign out_flat[209] = widths_cast_wrapper_out_flat[0];
  assign out_flat[111] = widths_cast_wrapper_out_flat[1];
  assign out_flat[343] = widths_cast_wrapper_out_flat[2];
  assign out_flat[327] = widths_cast_wrapper_out_flat[3];
  assign out_flat[282] = widths_cast_wrapper_out_flat[4];
  assign out_flat[393] = widths_cast_wrapper_out_flat[5];
  assign out_flat[405] = widths_cast_wrapper_out_flat[6];
  assign out_flat[240] = widths_cast_wrapper_out_flat[7];
  assign out_flat[133] = widths_cast_wrapper_out_flat[8];
  assign out_flat[101] = widths_cast_wrapper_out_flat[9];
  assign out_flat[331] = widths_cast_wrapper_out_flat[10];
  assign out_flat[151] = widths_cast_wrapper_out_flat[11];
  assign out_flat[404] = numbers_logical_op_wrapper_out_flat[0];
  assign out_flat[316] = numbers_logical_op_wrapper_out_flat[1];
  assign out_flat[5] = numbers_logical_op_wrapper_out_flat[2];
  assign out_flat[166] = widths_struct_mod_wrapper_out_flat[0];
  assign out_flat[409] = widths_struct_mod_wrapper_out_flat[1];
  assign out_flat[132] = widths_struct_mod_wrapper_out_flat[2];
  assign out_flat[91] = widths_struct_mod_wrapper_out_flat[3];
  assign out_flat[300] = widths_struct_mod_wrapper_out_flat[4];
  assign out_flat[177] = widths_struct_mod_wrapper_out_flat[5];
  assign out_flat[41] = widths_struct_mod_wrapper_out_flat[6];
  assign out_flat[73] = widths_struct_mod_wrapper_out_flat[7];
  assign out_flat[206] = widths_struct_mod_wrapper_out_flat[8];
  assign out_flat[342] = widths_struct_mod_wrapper_out_flat[9];
  assign out_flat[1] = widths_struct_mod_wrapper_out_flat[10];
  assign out_flat[397] = widths_struct_mod_wrapper_out_flat[11];
  assign out_flat[234] = widths_partselect_wrapper_out_flat[0];
  assign out_flat[381] = widths_partselect_wrapper_out_flat[1];
  assign out_flat[123] = widths_partselect_wrapper_out_flat[2];
  assign out_flat[269] = widths_partselect_wrapper_out_flat[3];
  assign out_flat[36] = widths_partselect_wrapper_out_flat[4];
  assign out_flat[145] = widths_partselect_wrapper_out_flat[5];
  assign out_flat[110] = widths_partselect_wrapper_out_flat[6];
  assign out_flat[328] = widths_partselect_wrapper_out_flat[7];
  assign out_flat[256] = widths_partselect_wrapper_out_flat[8];
  assign out_flat[440] = numbers_bitwise_reduce_wrapper_out_flat[0];
  assign out_flat[138] = numbers_bitwise_reduce_wrapper_out_flat[1];
  assign out_flat[278] = numbers_bitwise_reduce_wrapper_out_flat[2];
  assign out_flat[194] = numbers_arithmetic_reduce_wrapper_out_flat[0];
  assign out_flat[227] = numbers_arithmetic_reduce_wrapper_out_flat[1];
  assign out_flat[155] = numbers_arithmetic_reduce_wrapper_out_flat[2];
  assign out_flat[288] = numbers_arithmetic_reduce_wrapper_out_flat[3];
  assign out_flat[126] = numbers_arithmetic_reduce_wrapper_out_flat[4];
  assign out_flat[364] = numbers_arithmetic_reduce_wrapper_out_flat[5];
  assign out_flat[295] = numbers_arithmetic_reduce_wrapper_out_flat[6];
  assign out_flat[344] = numbers_arithmetic_reduce_wrapper_out_flat[7];
  assign out_flat[105] = numbers_arithmetic_reduce_wrapper_out_flat[8];
  assign out_flat[339] = numbers_arithmetic_reduce_wrapper_out_flat[9];
  assign out_flat[335] = widths_conditional_wrapper_out_flat[0];
  assign out_flat[172] = widths_conditional_wrapper_out_flat[1];
  assign out_flat[391] = widths_conditional_wrapper_out_flat[2];
  assign out_flat[362] = widths_conditional_wrapper_out_flat[3];
  assign out_flat[0] = const_arith_wrapper_out_flat[0];
  assign out_flat[158] = const_arith_wrapper_out_flat[1];
  assign out_flat[392] = const_arith_wrapper_out_flat[2];
  assign out_flat[461] = const_arith_wrapper_out_flat[3];
  assign out_flat[462] = const_arith_wrapper_out_flat[4];
  assign out_flat[12] = const_arith_wrapper_out_flat[5];
  assign out_flat[185] = const_arith_wrapper_out_flat[6];
  assign out_flat[413] = const_arith_wrapper_out_flat[7];
  assign out_flat[169] = const_arith_wrapper_out_flat[8];
  assign out_flat[410] = const_arith_wrapper_out_flat[9];
  assign out_flat[231] = const_arith_wrapper_out_flat[10];
  assign out_flat[396] = const_arith_wrapper_out_flat[11];
  assign out_flat[40] = const_arith_wrapper_out_flat[12];
  assign out_flat[375] = const_arith_wrapper_out_flat[13];
  assign out_flat[27] = const_arith_wrapper_out_flat[14];
  assign out_flat[154] = const_arith_wrapper_out_flat[15];
  assign out_flat[296] = const_arith_wrapper_out_flat[16];
  assign out_flat[225] = const_arith_wrapper_out_flat[17];
  assign out_flat[354] = const_arith_wrapper_out_flat[18];
  assign out_flat[457] = const_arith_wrapper_out_flat[19];
  assign out_flat[178] = const_arith_wrapper_out_flat[20];
  assign out_flat[243] = const_arith_wrapper_out_flat[21];
  assign out_flat[437] = const_arith_wrapper_out_flat[22];
  assign out_flat[330] = const_arith_wrapper_out_flat[23];
  assign out_flat[92] = const_arith_wrapper_out_flat[24];
  assign out_flat[108] = const_arith_wrapper_out_flat[25];
  assign out_flat[347] = const_arith_wrapper_out_flat[26];
  assign out_flat[63] = const_arith_wrapper_out_flat[27];
  assign out_flat[184] = const_arith_wrapper_out_flat[28];
  assign out_flat[49] = const_arith_wrapper_out_flat[29];
  assign out_flat[58] = const_arith_wrapper_out_flat[30];
  assign out_flat[356] = const_arith_wrapper_out_flat[31];
  assign out_flat[367] = const_arith_wrapper_out_flat[32];
  assign out_flat[459] = const_arith_wrapper_out_flat[33];
  assign out_flat[75] = const_arith_wrapper_out_flat[34];
  assign out_flat[51] = const_arith_wrapper_out_flat[35];
  assign out_flat[53] = const_arith_wrapper_out_flat[36];
  assign out_flat[134] = const_arith_wrapper_out_flat[37];
  assign out_flat[218] = const_arith_wrapper_out_flat[38];
  assign out_flat[193] = const_arith_wrapper_out_flat[39];
  assign out_flat[214] = widths_union_mod_wrapper_out_flat[0];
  assign out_flat[17] = widths_union_mod_wrapper_out_flat[1];
  assign out_flat[249] = widths_union_mod_wrapper_out_flat[2];
  assign out_flat[299] = widths_union_mod_wrapper_out_flat[3];
  assign out_flat[399] = widths_union_mod_wrapper_out_flat[4];
  assign out_flat[142] = widths_union_mod_wrapper_out_flat[5];
  assign out_flat[372] = widths_union_mod_wrapper_out_flat[6];
  assign out_flat[407] = widths_union_mod_wrapper_out_flat[7];
  assign out_flat[181] = widths_union_mod_wrapper_out_flat[8];
  assign out_flat[374] = widths_union_mod_wrapper_out_flat[9];
  assign out_flat[205] = widths_union_mod_wrapper_out_flat[10];
  assign out_flat[203] = widths_union_mod_wrapper_out_flat[11];
  assign out_flat[162] = widths_union_mod_wrapper_out_flat[12];
  assign out_flat[78] = widths_union_mod_wrapper_out_flat[13];
  assign out_flat[447] = widths_union_mod_wrapper_out_flat[14];
  assign out_flat[201] = widths_union_mod_wrapper_out_flat[15];
  assign out_flat[387] = const_shift_wrapper_out_flat[0];
  assign out_flat[274] = const_shift_wrapper_out_flat[1];
  assign out_flat[247] = const_shift_wrapper_out_flat[2];
  assign out_flat[104] = const_shift_wrapper_out_flat[3];
  assign out_flat[400] = const_shift_wrapper_out_flat[4];
  assign out_flat[329] = const_shift_wrapper_out_flat[5];
  assign out_flat[25] = const_shift_wrapper_out_flat[6];
  assign out_flat[304] = const_shift_wrapper_out_flat[7];
  assign out_flat[352] = const_shift_wrapper_out_flat[8];
  assign out_flat[46] = const_shift_wrapper_out_flat[9];
  assign out_flat[208] = const_shift_wrapper_out_flat[10];
  assign out_flat[386] = const_shift_wrapper_out_flat[11];
  assign out_flat[37] = const_shift_wrapper_out_flat[12];
  assign out_flat[237] = const_shift_wrapper_out_flat[13];
  assign out_flat[258] = const_shift_wrapper_out_flat[14];
  assign out_flat[100] = const_shift_wrapper_out_flat[15];
  assign out_flat[26] = const_shift_wrapper_out_flat[16];
  assign out_flat[290] = const_shift_wrapper_out_flat[17];
  assign out_flat[469] = const_shift_wrapper_out_flat[18];
  assign out_flat[238] = const_shift_wrapper_out_flat[19];
  assign out_flat[379] = const_shift_wrapper_out_flat[20];
  assign out_flat[232] = const_shift_wrapper_out_flat[21];
  assign out_flat[348] = const_shift_wrapper_out_flat[22];
  assign out_flat[72] = const_shift_wrapper_out_flat[23];
  assign out_flat[117] = widths_logic_mod_wrapper_out_flat[0];
  assign out_flat[384] = widths_logic_mod_wrapper_out_flat[1];
  assign out_flat[248] = widths_logic_mod_wrapper_out_flat[2];
  assign out_flat[202] = widths_logic_mod_wrapper_out_flat[3];
  assign out_flat[244] = widths_logic_mod_wrapper_out_flat[4];
  assign out_flat[349] = widths_logic_mod_wrapper_out_flat[5];
  assign out_flat[418] = widths_array_wrapper_out_flat[0];
  assign out_flat[34] = widths_array_wrapper_out_flat[1];
  assign out_flat[211] = widths_array_wrapper_out_flat[2];
  assign out_flat[353] = widths_array_wrapper_out_flat[3];
  assign out_flat[161] = widths_array_wrapper_out_flat[4];
  assign out_flat[222] = widths_array_wrapper_out_flat[5];
  assign out_flat[377] = widths_array_wrapper_out_flat[6];
  assign out_flat[52] = widths_array_wrapper_out_flat[7];
  assign out_flat[424] = widths_array_wrapper_out_flat[8];
  assign out_flat[260] = widths_array_wrapper_out_flat[9];
  assign out_flat[261] = widths_array_wrapper_out_flat[10];
  assign out_flat[449] = widths_array_wrapper_out_flat[11];
  assign out_flat[254] = widths_array_wrapper_out_flat[12];
  assign out_flat[426] = widths_array_wrapper_out_flat[13];
  assign out_flat[106] = widths_array_wrapper_out_flat[14];
  assign out_flat[186] = widths_array_wrapper_out_flat[15];
  assign out_flat[175] = numbers_select_wrapper_out_flat[0];
  assign out_flat[433] = numbers_select_wrapper_out_flat[1];
  assign out_flat[11] = numbers_select_wrapper_out_flat[2];
  assign out_flat[345] = numbers_select_wrapper_out_flat[3];
  assign out_flat[474] = numbers_select_wrapper_out_flat[4];
  assign out_flat[332] = numbers_select_wrapper_out_flat[5];
  assign out_flat[6] = numbers_select_wrapper_out_flat[6];
  assign out_flat[287] = numbers_select_wrapper_out_flat[7];
  assign out_flat[192] = numbers_select_wrapper_out_flat[8];
  assign out_flat[94] = widths_arith_wrapper_out_flat[0];
  assign out_flat[65] = const_nested_wrapper_out_flat[0];
  assign out_flat[442] = const_nested_wrapper_out_flat[1];
  assign out_flat[378] = const_nested_wrapper_out_flat[2];
  assign out_flat[246] = const_nested_wrapper_out_flat[3];
  assign out_flat[86] = const_nested_wrapper_out_flat[4];
  assign out_flat[120] = const_nested_wrapper_out_flat[5];
  assign out_flat[21] = const_nested_wrapper_out_flat[6];
  assign out_flat[146] = const_nested_wrapper_out_flat[7];
  assign out_flat[365] = numbers_numbers_arithmetic_wrapper_out_flat[0];
  assign out_flat[187] = numbers_numbers_arithmetic_wrapper_out_flat[1];
  assign out_flat[351] = numbers_numbers_arithmetic_wrapper_out_flat[2];
  assign out_flat[15] = numbers_numbers_arithmetic_wrapper_out_flat[3];
  assign out_flat[453] = numbers_numbers_arithmetic_wrapper_out_flat[4];
  assign out_flat[285] = numbers_numbers_arithmetic_wrapper_out_flat[5];
  assign out_flat[320] = numbers_numbers_arithmetic_wrapper_out_flat[6];
  assign out_flat[118] = numbers_numbers_arithmetic_wrapper_out_flat[7];
  assign out_flat[428] = numbers_numbers_arithmetic_wrapper_out_flat[8];
  assign out_flat[14] = numbers_numbers_arithmetic_wrapper_out_flat[9];
  assign out_flat[44] = numbers_numbers_arithmetic_wrapper_out_flat[10];
  assign out_flat[197] = numbers_numbers_arithmetic_wrapper_out_flat[11];
  assign out_flat[376] = numbers_numbers_arithmetic_wrapper_out_flat[12];
  assign out_flat[62] = numbers_numbers_arithmetic_wrapper_out_flat[13];
  assign out_flat[323] = numbers_numbers_arithmetic_wrapper_out_flat[14];
  assign out_flat[436] = numbers_numbers_arithmetic_wrapper_out_flat[15];
  assign out_flat[337] = numbers_numbers_arithmetic_wrapper_out_flat[16];
  assign out_flat[236] = numbers_numbers_arithmetic_wrapper_out_flat[17];
  assign out_flat[85] = numbers_numbers_arithmetic_wrapper_out_flat[18];
  assign out_flat[310] = numbers_numbers_arithmetic_wrapper_out_flat[19];
  assign out_flat[228] = numbers_numbers_arithmetic_wrapper_out_flat[20];
  assign out_flat[56] = numbers_numbers_arithmetic_wrapper_out_flat[21];
  assign out_flat[170] = numbers_numbers_arithmetic_wrapper_out_flat[22];
  assign out_flat[144] = numbers_numbers_arithmetic_wrapper_out_flat[23];
  assign out_flat[165] = numbers_numbers_arithmetic_wrapper_out_flat[24];
  assign out_flat[79] = numbers_bitwise_logic_wrapper_out_flat[0];
  assign out_flat[283] = numbers_bitwise_logic_wrapper_out_flat[1];
  assign out_flat[97] = numbers_bitwise_logic_wrapper_out_flat[2];
  assign out_flat[402] = numbers_bitwise_logic_wrapper_out_flat[3];
  assign out_flat[385] = numbers_bitwise_logic_wrapper_out_flat[4];
  assign out_flat[180] = numbers_bitwise_logic_wrapper_out_flat[5];
  assign out_flat[417] = numbers_bitwise_logic_wrapper_out_flat[6];
  assign out_flat[47] = numbers_bitwise_logic_wrapper_out_flat[7];
  assign out_flat[235] = numbers_bitwise_logic_wrapper_out_flat[8];
  assign out_flat[196] = numbers_bitwise_logic_wrapper_out_flat[9];
  assign out_flat[242] = numbers_bitwise_logic_wrapper_out_flat[10];
  assign out_flat[220] = numbers_bitwise_logic_wrapper_out_flat[11];
  assign out_flat[471] = numbers_bitwise_logic_wrapper_out_flat[12];
  assign out_flat[96] = numbers_bitwise_logic_wrapper_out_flat[13];
  assign out_flat[382] = numbers_bitwise_logic_wrapper_out_flat[14];
  assign out_flat[239] = numbers_bitwise_logic_wrapper_out_flat[15];
  assign out_flat[333] = numbers_bitwise_logic_wrapper_out_flat[16];
  assign out_flat[18] = numbers_bitwise_logic_wrapper_out_flat[17];
  assign out_flat[434] = numbers_bitwise_logic_wrapper_out_flat[18];
  assign out_flat[280] = numbers_bitwise_logic_wrapper_out_flat[19];
  assign out_flat[427] = numbers_bitwise_logic_wrapper_out_flat[20];
  assign out_flat[90] = numbers_bitwise_logic_wrapper_out_flat[21];
  assign out_flat[473] = numbers_bitwise_logic_wrapper_out_flat[22];
  assign out_flat[216] = numbers_bitwise_logic_wrapper_out_flat[23];
  assign out_flat[114] = widths_concat_repl_wrapper_out_flat[0];
  assign out_flat[99] = widths_concat_repl_wrapper_out_flat[1];
  assign out_flat[383] = widths_concat_repl_wrapper_out_flat[2];
  assign out_flat[23] = widths_concat_repl_wrapper_out_flat[3];
  assign out_flat[31] = widths_concat_repl_wrapper_out_flat[4];
  assign out_flat[460] = widths_concat_repl_wrapper_out_flat[5];
  assign out_flat[22] = widths_concat_repl_wrapper_out_flat[6];
  assign out_flat[29] = widths_concat_repl_wrapper_out_flat[7];
  assign out_flat[2] = widths_concat_repl_wrapper_out_flat[8];
  assign out_flat[371] = widths_concat_repl_wrapper_out_flat[9];
  assign out_flat[441] = widths_concat_repl_wrapper_out_flat[10];
  assign out_flat[452] = widths_concat_repl_wrapper_out_flat[11];
  assign out_flat[251] = widths_concat_repl_wrapper_out_flat[12];
  assign out_flat[439] = widths_concat_repl_wrapper_out_flat[13];
  assign out_flat[476] = widths_concat_repl_wrapper_out_flat[14];
  assign out_flat[204] = widths_concat_repl_wrapper_out_flat[15];
  assign out_flat[267] = widths_concat_repl_wrapper_out_flat[16];
  assign out_flat[301] = widths_concat_repl_wrapper_out_flat[17];
  assign out_flat[59] = const_partselect_wrapper_out_flat[0];
  assign out_flat[159] = const_partselect_wrapper_out_flat[1];
  assign out_flat[294] = const_partselect_wrapper_out_flat[2];
  assign out_flat[319] = const_partselect_wrapper_out_flat[3];
  assign out_flat[124] = const_partselect_wrapper_out_flat[4];
  assign out_flat[422] = const_partselect_wrapper_out_flat[5];
  assign out_flat[456] = const_partselect_wrapper_out_flat[6];
  assign out_flat[67] = const_partselect_wrapper_out_flat[7];
  assign out_flat[152] = numbers_constant_wrapper_out_flat[0];
  assign out_flat[312] = numbers_constant_wrapper_out_flat[1];
  assign out_flat[10] = numbers_constant_wrapper_out_flat[2];
  assign out_flat[412] = numbers_constant_wrapper_out_flat[3];
  assign out_flat[408] = numbers_constant_wrapper_out_flat[4];
  assign out_flat[54] = numbers_constant_wrapper_out_flat[5];
  assign out_flat[43] = numbers_constant_wrapper_out_flat[6];
  assign out_flat[116] = numbers_constant_wrapper_out_flat[7];
  assign out_flat[167] = numbers_constant_wrapper_out_flat[8];
  assign out_flat[438] = numbers_constant_wrapper_out_flat[9];
  assign out_flat[281] = numbers_constant_wrapper_out_flat[10];
  assign out_flat[149] = numbers_constant_wrapper_out_flat[11];
  assign out_flat[311] = numbers_constant_wrapper_out_flat[12];
  assign out_flat[432] = numbers_constant_wrapper_out_flat[13];
  assign out_flat[259] = numbers_constant_wrapper_out_flat[14];
  assign out_flat[109] = numbers_constant_wrapper_out_flat[15];
  assign out_flat[135] = numbers_constant_wrapper_out_flat[16];
  assign out_flat[450] = numbers_constant_wrapper_out_flat[17];
  assign out_flat[465] = numbers_constant_wrapper_out_flat[18];
  assign out_flat[125] = numbers_constant_wrapper_out_flat[19];
  assign out_flat[262] = numbers_constant_wrapper_out_flat[20];
  assign out_flat[411] = numbers_constant_wrapper_out_flat[21];
  assign out_flat[24] = numbers_constant_wrapper_out_flat[22];
  assign out_flat[20] = numbers_constant_wrapper_out_flat[23];
  assign out_flat[74] = numbers_constant_wrapper_out_flat[24];
  assign out_flat[466] = numbers_constant_wrapper_out_flat[25];
  assign out_flat[263] = numbers_constant_wrapper_out_flat[26];
  assign out_flat[150] = numbers_constant_wrapper_out_flat[27];
  assign out_flat[268] = numbers_constant_wrapper_out_flat[28];
  assign out_flat[416] = numbers_constant_wrapper_out_flat[29];
  assign out_flat[279] = numbers_constant_wrapper_out_flat[30];
  assign out_flat[122] = numbers_constant_wrapper_out_flat[31];
  assign out_flat[147] = numbers_constant_wrapper_out_flat[32];
  assign out_flat[84] = numbers_constant_wrapper_out_flat[33];
  assign out_flat[171] = numbers_constant_wrapper_out_flat[34];
  assign out_flat[419] = numbers_constant_wrapper_out_flat[35];
  assign out_flat[467] = numbers_constant_wrapper_out_flat[36];
  assign out_flat[215] = numbers_constant_wrapper_out_flat[37];
  assign out_flat[390] = numbers_constant_wrapper_out_flat[38];
  assign out_flat[334] = numbers_constant_wrapper_out_flat[39];
  assign out_flat[250] = numbers_constant_wrapper_out_flat[40];
  assign out_flat[420] = numbers_constant_wrapper_out_flat[41];
  assign out_flat[128] = numbers_constant_wrapper_out_flat[42];
  assign out_flat[207] = numbers_constant_wrapper_out_flat[43];
  assign out_flat[39] = numbers_constant_wrapper_out_flat[44];
  assign out_flat[121] = numbers_constant_wrapper_out_flat[45];
  assign out_flat[270] = numbers_constant_wrapper_out_flat[46];
  assign out_flat[219] = numbers_constant_wrapper_out_flat[47];
  assign out_flat[265] = numbers_constant_wrapper_out_flat[48];
  assign out_flat[137] = numbers_constant_wrapper_out_flat[49];
  assign out_flat[42] = numbers_constant_wrapper_out_flat[50];
  assign out_flat[163] = numbers_constant_wrapper_out_flat[51];
  assign out_flat[289] = numbers_constant_wrapper_out_flat[52];
  assign out_flat[463] = numbers_constant_wrapper_out_flat[53];
  assign out_flat[68] = numbers_constant_wrapper_out_flat[54];
  assign out_flat[95] = numbers_constant_wrapper_out_flat[55];
  assign out_flat[160] = numbers_constant_wrapper_out_flat[56];
  assign out_flat[153] = numbers_constant_wrapper_out_flat[57];
  assign out_flat[359] = numbers_constant_wrapper_out_flat[58];
  assign out_flat[446] = numbers_constant_wrapper_out_flat[59];
  assign out_flat[191] = numbers_constant_wrapper_out_flat[60];
  assign out_flat[3] = numbers_constant_wrapper_out_flat[61];
  assign out_flat[13] = numbers_constant_wrapper_out_flat[62];
  assign out_flat[350] = numbers_constant_wrapper_out_flat[63];
  assign out_flat[143] = numbers_constant_wrapper_out_flat[64];
  assign out_flat[28] = numbers_constant_wrapper_out_flat[65];
  assign out_flat[293] = numbers_constant_wrapper_out_flat[66];
  assign out_flat[8] = numbers_constant_wrapper_out_flat[67];
  assign out_flat[50] = numbers_constant_wrapper_out_flat[68];
  assign out_flat[398] = numbers_constant_wrapper_out_flat[69];
  assign out_flat[176] = numbers_constant_wrapper_out_flat[70];
  assign out_flat[313] = numbers_constant_wrapper_out_flat[71];
  assign out_flat[210] = numbers_constant_wrapper_out_flat[72];
  assign out_flat[64] = numbers_constant_wrapper_out_flat[73];
  assign out_flat[338] = numbers_constant_wrapper_out_flat[74];
  assign out_flat[273] = numbers_constant_wrapper_out_flat[75];
  assign out_flat[182] = numbers_constant_wrapper_out_flat[76];
  assign out_flat[445] = numbers_constant_wrapper_out_flat[77];
  assign out_flat[80] = numbers_constant_wrapper_out_flat[78];
  assign out_flat[430] = numbers_constant_wrapper_out_flat[79];
  assign out_flat[136] = const_compare_wrapper_out_flat[0];
  assign out_flat[9] = const_compare_wrapper_out_flat[1];
  assign out_flat[468] = const_compare_wrapper_out_flat[2];
  assign out_flat[388] = const_compare_wrapper_out_flat[3];
  assign out_flat[253] = const_compare_wrapper_out_flat[4];
  assign out_flat[212] = const_compare_wrapper_out_flat[5];
  assign out_flat[32] = const_compare_wrapper_out_flat[6];
  assign out_flat[255] = const_compare_wrapper_out_flat[7];
  assign out_flat[174] = widths_param_wrapper_out_flat[0];
  assign out_flat[317] = const_reduce_wrapper_out_flat[0];
  assign out_flat[107] = const_reduce_wrapper_out_flat[1];
  assign out_flat[77] = const_reduce_wrapper_out_flat[2];
  assign out_flat[38] = const_reduce_wrapper_out_flat[3];
  assign out_flat[61] = const_reduce_wrapper_out_flat[4];
  assign out_flat[355] = const_reduce_wrapper_out_flat[5];
  assign out_flat[245] = const_concat_repl_wrapper_out_flat[0];
  assign out_flat[148] = const_concat_repl_wrapper_out_flat[1];
  assign out_flat[464] = const_concat_repl_wrapper_out_flat[2];
  assign out_flat[322] = const_concat_repl_wrapper_out_flat[3];
  assign out_flat[7] = const_concat_repl_wrapper_out_flat[4];
  assign out_flat[373] = const_concat_repl_wrapper_out_flat[5];
  assign out_flat[131] = const_concat_repl_wrapper_out_flat[6];
  assign out_flat[35] = const_concat_repl_wrapper_out_flat[7];
  assign out_flat[341] = const_concat_repl_wrapper_out_flat[8];
  assign out_flat[127] = const_concat_repl_wrapper_out_flat[9];
  assign out_flat[284] = const_concat_repl_wrapper_out_flat[10];
  assign out_flat[291] = const_concat_repl_wrapper_out_flat[11];
  assign out_flat[340] = const_concat_repl_wrapper_out_flat[12];
  assign out_flat[157] = const_concat_repl_wrapper_out_flat[13];
  assign out_flat[455] = const_concat_repl_wrapper_out_flat[14];
  assign out_flat[102] = const_concat_repl_wrapper_out_flat[15];
  assign out_flat[98] = const_concat_repl_wrapper_out_flat[16];
  assign out_flat[83] = const_concat_repl_wrapper_out_flat[17];
  assign out_flat[57] = const_concat_repl_wrapper_out_flat[18];
  assign out_flat[82] = const_concat_repl_wrapper_out_flat[19];
  assign out_flat[277] = const_concat_repl_wrapper_out_flat[20];
  assign out_flat[271] = const_concat_repl_wrapper_out_flat[21];
  assign out_flat[119] = numbers_reduce_case_wrapper_out_flat[0];
  assign out_flat[156] = numbers_reduce_case_wrapper_out_flat[1];
  assign out_flat[129] = widths_enum_mod_wrapper_out_flat[0];
  assign out_flat[475] = widths_enum_mod_wrapper_out_flat[1];
  assign out_flat[429] = widths_enum_mod_wrapper_out_flat[2];
  assign out_flat[346] = widths_enum_mod_wrapper_out_flat[3];
  assign out_flat[325] = widths_enum_mod_wrapper_out_flat[4];
  assign out_flat[318] = const_conditional_wrapper_out_flat[0];
  assign out_flat[93] = const_conditional_wrapper_out_flat[1];
  assign out_flat[275] = const_conditional_wrapper_out_flat[2];
  assign out_flat[326] = const_conditional_wrapper_out_flat[3];
  assign out_flat[360] = const_conditional_wrapper_out_flat[4];
  assign out_flat[264] = const_conditional_wrapper_out_flat[5];
  assign out_flat[199] = const_conditional_wrapper_out_flat[6];
  assign out_flat[173] = const_conditional_wrapper_out_flat[7];
  assign out_flat[76] = const_conditional_wrapper_out_flat[8];
  assign out_flat[297] = const_conditional_wrapper_out_flat[9];
  assign out_flat[16] = const_conditional_wrapper_out_flat[10];
  assign out_flat[190] = const_conditional_wrapper_out_flat[11];
  assign out_flat[321] = const_conditional_wrapper_out_flat[12];
  assign out_flat[112] = const_conditional_wrapper_out_flat[13];
  assign out_flat[309] = const_conditional_wrapper_out_flat[14];
  assign out_flat[198] = const_conditional_wrapper_out_flat[15];
  assign out_flat[308] = const_conditional_wrapper_out_flat[16];
  assign out_flat[315] = const_conditional_wrapper_out_flat[17];
  assign out_flat[141] = const_conditional_wrapper_out_flat[18];
  assign out_flat[200] = const_conditional_wrapper_out_flat[19];
  assign out_flat[217] = const_conditional_wrapper_out_flat[20];
  assign out_flat[394] = const_conditional_wrapper_out_flat[21];
  assign out_flat[448] = const_conditional_wrapper_out_flat[22];
  assign out_flat[307] = const_conditional_wrapper_out_flat[23];
  assign out_flat[358] = numbers_shift_wrapper_out_flat[0];
  assign out_flat[87] = numbers_shift_wrapper_out_flat[1];
  assign out_flat[454] = numbers_shift_wrapper_out_flat[2];
  assign out_flat[451] = numbers_shift_wrapper_out_flat[3];
  assign out_flat[179] = numbers_shift_wrapper_out_flat[4];
  assign out_flat[431] = numbers_shift_wrapper_out_flat[5];
  assign out_flat[303] = numbers_shift_wrapper_out_flat[6];
  assign out_flat[4] = numbers_shift_wrapper_out_flat[7];
  assign out_flat[425] = numbers_shift_wrapper_out_flat[8];
  assign out_flat[213] = numbers_shift_wrapper_out_flat[9];
  assign out_flat[389] = numbers_shift_wrapper_out_flat[10];
  assign out_flat[415] = numbers_shift_wrapper_out_flat[11];
  assign out_flat[188] = numbers_shift_wrapper_out_flat[12];
  assign out_flat[30] = numbers_shift_wrapper_out_flat[13];
  assign out_flat[302] = numbers_shift_wrapper_out_flat[14];
  assign out_flat[395] = numbers_shift_wrapper_out_flat[15];
  assign out_flat[230] = const_logic_wrapper_out_flat[0];
  assign out_flat[292] = const_logic_wrapper_out_flat[1];
  assign out_flat[241] = const_logic_wrapper_out_flat[2];
  assign out_flat[140] = const_logic_wrapper_out_flat[3];
  assign out_flat[226] = const_logic_wrapper_out_flat[4];
  assign out_flat[45] = const_logic_wrapper_out_flat[5];
  assign out_flat[472] = const_logic_wrapper_out_flat[6];
  assign out_flat[229] = const_logic_wrapper_out_flat[7];
  assign out_flat[305] = const_logic_wrapper_out_flat[8];
  assign out_flat[286] = const_logic_wrapper_out_flat[9];
  assign out_flat[414] = const_logic_wrapper_out_flat[10];
  assign out_flat[103] = const_logic_wrapper_out_flat[11];
  assign out_flat[33] = const_logic_wrapper_out_flat[12];
  assign out_flat[272] = const_logic_wrapper_out_flat[13];
  assign out_flat[361] = const_logic_wrapper_out_flat[14];
  assign out_flat[88] = const_logic_wrapper_out_flat[15];
  assign out_flat[221] = const_logic_wrapper_out_flat[16];
  assign out_flat[130] = const_logic_wrapper_out_flat[17];
  assign out_flat[139] = const_logic_wrapper_out_flat[18];
  assign out_flat[444] = widths_shift_wrapper_out_flat[0];
  assign out_flat[369] = widths_shift_wrapper_out_flat[1];
  assign out_flat[314] = widths_shift_wrapper_out_flat[2];
  assign out_flat[223] = widths_shift_wrapper_out_flat[3];
  assign out_flat[421] = widths_shift_wrapper_out_flat[4];
  assign out_flat[60] = widths_shift_wrapper_out_flat[5];
  assign out_flat[115] = widths_shift_wrapper_out_flat[6];
  assign out_flat[195] = widths_shift_wrapper_out_flat[7];
  assign out_flat[370] = widths_shift_wrapper_out_flat[8];
  assign out_flat[113] = widths_shift_wrapper_out_flat[9];
  assign out_flat[257] = widths_shift_wrapper_out_flat[10];
  assign out_flat[189] = widths_shift_wrapper_out_flat[11];
  assign out_flat[324] = widths_shift_wrapper_out_flat[12];
  assign out_flat[357] = widths_shift_wrapper_out_flat[13];
  assign out_flat[48] = widths_shift_wrapper_out_flat[14];
  assign out_flat[55] = widths_shift_wrapper_out_flat[15];

  // Instantiate each module's wrapper
  const_arith_wrapper u_const_arith_wrapper (
    .in_flat  (const_arith_wrapper_in_flat),
    .out_flat (const_arith_wrapper_out_flat)
  );
  const_compare_wrapper u_const_compare_wrapper (
    .in_flat  (const_compare_wrapper_in_flat),
    .out_flat (const_compare_wrapper_out_flat)
  );
  const_concat_repl_wrapper u_const_concat_repl_wrapper (
    .in_flat  (const_concat_repl_wrapper_in_flat),
    .out_flat (const_concat_repl_wrapper_out_flat)
  );
  const_conditional_wrapper u_const_conditional_wrapper (
    .in_flat  (const_conditional_wrapper_in_flat),
    .out_flat (const_conditional_wrapper_out_flat)
  );
  const_logic_wrapper u_const_logic_wrapper (
    .in_flat  (const_logic_wrapper_in_flat),
    .out_flat (const_logic_wrapper_out_flat)
  );
  const_nested_wrapper u_const_nested_wrapper (
    .in_flat  (const_nested_wrapper_in_flat),
    .out_flat (const_nested_wrapper_out_flat)
  );
  const_partselect_wrapper u_const_partselect_wrapper (
    .in_flat  (const_partselect_wrapper_in_flat),
    .out_flat (const_partselect_wrapper_out_flat)
  );
  const_reduce_wrapper u_const_reduce_wrapper (
    .in_flat  (const_reduce_wrapper_in_flat),
    .out_flat (const_reduce_wrapper_out_flat)
  );
  const_shift_wrapper u_const_shift_wrapper (
    .in_flat  (const_shift_wrapper_in_flat),
    .out_flat (const_shift_wrapper_out_flat)
  );
  numbers_arithmetic_reduce_wrapper u_numbers_arithmetic_reduce_wrapper (
    .in_flat  (numbers_arithmetic_reduce_wrapper_in_flat),
    .out_flat (numbers_arithmetic_reduce_wrapper_out_flat)
  );
  numbers_bitwise_logic_wrapper u_numbers_bitwise_logic_wrapper (
    .in_flat  (numbers_bitwise_logic_wrapper_in_flat),
    .out_flat (numbers_bitwise_logic_wrapper_out_flat)
  );
  numbers_bitwise_reduce_wrapper u_numbers_bitwise_reduce_wrapper (
    .in_flat  (numbers_bitwise_reduce_wrapper_in_flat),
    .out_flat (numbers_bitwise_reduce_wrapper_out_flat)
  );
  numbers_concat_repl_wrapper u_numbers_concat_repl_wrapper (
    .in_flat  (numbers_concat_repl_wrapper_in_flat),
    .out_flat (numbers_concat_repl_wrapper_out_flat)
  );
  numbers_constant_wrapper u_numbers_constant_wrapper (
    .in_flat  (numbers_constant_wrapper_in_flat),
    .out_flat (numbers_constant_wrapper_out_flat)
  );
  numbers_logical_op_wrapper u_numbers_logical_op_wrapper (
    .in_flat  (numbers_logical_op_wrapper_in_flat),
    .out_flat (numbers_logical_op_wrapper_out_flat)
  );
  numbers_numbers_arithmetic_wrapper u_numbers_numbers_arithmetic_wrapper (
    .in_flat  (numbers_numbers_arithmetic_wrapper_in_flat),
    .out_flat (numbers_numbers_arithmetic_wrapper_out_flat)
  );
  numbers_reduce_case_wrapper u_numbers_reduce_case_wrapper (
    .in_flat  (numbers_reduce_case_wrapper_in_flat),
    .out_flat (numbers_reduce_case_wrapper_out_flat)
  );
  numbers_relational_wrapper u_numbers_relational_wrapper (
    .in_flat  (numbers_relational_wrapper_in_flat),
    .out_flat (numbers_relational_wrapper_out_flat)
  );
  numbers_select_wrapper u_numbers_select_wrapper (
    .in_flat  (numbers_select_wrapper_in_flat),
    .out_flat (numbers_select_wrapper_out_flat)
  );
  numbers_shift_wrapper u_numbers_shift_wrapper (
    .in_flat  (numbers_shift_wrapper_in_flat),
    .out_flat (numbers_shift_wrapper_out_flat)
  );
  widths_arith_wrapper u_widths_arith_wrapper (
    .in_flat  (widths_arith_wrapper_in_flat),
    .out_flat (widths_arith_wrapper_out_flat)
  );
  widths_array_wrapper u_widths_array_wrapper (
    .in_flat  (widths_array_wrapper_in_flat),
    .out_flat (widths_array_wrapper_out_flat)
  );
  widths_cast_wrapper u_widths_cast_wrapper (
    .in_flat  (widths_cast_wrapper_in_flat),
    .out_flat (widths_cast_wrapper_out_flat)
  );
  widths_concat_repl_wrapper u_widths_concat_repl_wrapper (
    .in_flat  (widths_concat_repl_wrapper_in_flat),
    .out_flat (widths_concat_repl_wrapper_out_flat)
  );
  widths_conditional_wrapper u_widths_conditional_wrapper (
    .in_flat  (widths_conditional_wrapper_in_flat),
    .out_flat (widths_conditional_wrapper_out_flat)
  );
  widths_enum_mod_wrapper u_widths_enum_mod_wrapper (
    .in_flat  (widths_enum_mod_wrapper_in_flat),
    .out_flat (widths_enum_mod_wrapper_out_flat)
  );
  widths_logic_mod_wrapper u_widths_logic_mod_wrapper (
    .in_flat  (widths_logic_mod_wrapper_in_flat),
    .out_flat (widths_logic_mod_wrapper_out_flat)
  );
  widths_param_wrapper u_widths_param_wrapper (
    .in_flat  (widths_param_wrapper_in_flat),
    .out_flat (widths_param_wrapper_out_flat)
  );
  widths_partselect_wrapper u_widths_partselect_wrapper (
    .in_flat  (widths_partselect_wrapper_in_flat),
    .out_flat (widths_partselect_wrapper_out_flat)
  );
  widths_shift_wrapper u_widths_shift_wrapper (
    .in_flat  (widths_shift_wrapper_in_flat),
    .out_flat (widths_shift_wrapper_out_flat)
  );
  widths_struct_mod_wrapper u_widths_struct_mod_wrapper (
    .in_flat  (widths_struct_mod_wrapper_in_flat),
    .out_flat (widths_struct_mod_wrapper_out_flat)
  );
  widths_union_mod_wrapper u_widths_union_mod_wrapper (
    .in_flat  (widths_union_mod_wrapper_in_flat),
    .out_flat (widths_union_mod_wrapper_out_flat)
  );

endmodule